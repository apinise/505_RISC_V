//////////////////////////////////////////////////////////////// 
// Engineer: Evan Apinis
// 
// Module Name: ctrl_logic.sv
// Project Name: RV32I 
// Description: 
// 
// Control logic for RV32I to decode instructions and control
// datapathing.
//
// Revision 0.01 - File Created
// 
////////////////////////////////////////////////////////////////

module ctrl_logic (
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

endmodule