//////////////////////////////////////////////////////////////// 
// Engineer: Evan Apinis
// 
// Module Name: proc_top.sv
// Project Name: RV32I 
// Description: 
// 
// RV32I processor top file including hart datapath and
// memory modules
//
// Revision 0.01 - File Created
// 
////////////////////////////////////////////////////////////////

module proc_top #(
  parameter DWIDTH = 32;
)(
  input logic Clk_Core,
  input logic Rst_Core_N
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

instruct_mem #(
  .DWIDTH(DWIDTH)
  .MEM_SIZE(16384)
)
instruct_mem (
  .Clk_Core(Clk_Core),
  .Rst_Core_N(Rst_Core_N),
  .Program_Count(),
  .Instruction()
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

endmodule