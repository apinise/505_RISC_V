module proc_top_r_tb (
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic clk;
logic rst_core_n;

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

proc_top #(
  .DWIDTH(32)
)
dut (
  .Clk_Core(clk)
  //.Rst_Core_N(rst_core_n)
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

initial begin
  clk = 0;
  rst_core_n = 0;
  # 10;
  rst_core_n = 1;
end

always begin
  #5;
  clk <= ~clk;
end

/*
initial begin
  wait (rst_core_n);
end
*/

endmodule