//////////////////////////////////////////////////////////////// 
// Engineer: Evan Apinis
// 
// Module Name: proc_top.sv
// Project Name: RV32I 
// Description: 
// 
// RV32I processor top file including hart datapath and
// memory modules
//
// Revision 0.01 - File Created
// 
////////////////////////////////////////////////////////////////

module proc_top #(
  parameter DWIDTH = 32
)(
  input logic Clk_Core,
  input logic Rst_Core_N
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic [DWIDTH-1:0]  program_count;
logic [31:0]        instruction;

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

core #(
  .DWIDTH()
)
core_1 (
  .Clk_Core(Clk_Core),
  .Rst_Core_N(Rst_Core_N),
  .Instruction(instruction),
  .Program_Count(program_count)
);

instruct_mem #(
  .DWIDTH(DWIDTH),
  .MEM_SIZE(16384)
)
instruct_mem (
  .Clk_Core(Clk_Core),
  .Rst_Core_N(Rst_Core_N),
  .Program_Count(program_count),
  .Instruction(instruction)
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

endmodule